`include "bsg_comm_link.vh"

//
// 8/4/2016 MBT
//
//
//

module bsg_frame_io #(parameter num_channels_p=4
                      ,parameter channel_width_p=8
                      ,parameter gateway_p=0
                      ,parameter nodes_p=1

                      ,parameter bsg_comm_link_i_s_width_lp = `bsg_comm_link_channel_in_s_width (channel_width_p)
                      ,parameter bsg_comm_link_o_s_width_lp = `bsg_comm_link_channel_out_s_width(channel_width_p)

                      ,parameter bsg_fsb_in_s_width_lp      = `bsg_fsb_in_s_width (ring_width_lp)
                      ,parameter bsg_fsb_out_s_width_lp     = `bsg_fsb_out_s_width(ring_width_lp)
                      )
   (
    input core_clk_i
    , input async_reset_i
    , input io_master_clk_i

    // I/O (comm_link side)
    , input  [num_channels_p-1:0][bsg_comm_link_i_s_width_lp-1:0] bsg_comm_link_i
    , output [num_channels_p-1:0][bsg_comm_link_o_s_width_lp-1:0] bsg_comm_link_o

    // I/O (fsb side)
    , input  [nodes_p-1:0][bsg_fsb_in_s_width_lp -1:0] fsb_li
    , output [nodes_p-1:0][bsg_fsb_out_s_width_lp-1:0] fsb_lo

    // generated by master (FPGA) and sent to slave (ASIC); unused by slave
    , output reg im_slave_reset_tline_r_o

    // post-calibration reset signal synchronous to the core clock
    , output core_reset_o
    );

   // **************************************************************
   // *
   // * convert bsg_comm_link structs to bsg_comm_link native format
   // *
   // * fixme: eventually we will push channel grouping down
   // * into bsg_comm_link, but the module is currently in flux
   // *

   `declare_bsg_comm_link_channel_in_s(channel_width_p);
   `declare_bsg_comm_link_channel_out_s(channel_width_p);

   bsg_comm_link_channel_in_s  [num_channels_p-1:0] bsg_comm_link_i_cast;
   bsg_comm_link_channel_out_s [num_channels_p-1:0] bsg_comm_link_o_cast;

   assign bsg_comm_link_i_cast = bsg_comm_link_i;
   assign bsg_comm_link_o      = bsg_comm_link_o_cast;

   // in channel
   logic [num_channels_p-1:0]  io_clk_tline_li;
   logic [num_channels_p-1:0]  io_valid_tline_li;
   logic [channel_width_p-1:0] io_data_tline_li [num_channels_p-1:0];
   logic [num_channels_p-1:0]  io_token_clk_tline_lo;

   genvar i;

   // input channel conversion
   for (i = 0; i < num_channels_p; i=i+1)
     begin:
        assign io_clk_tline_i      [i]                       = bsg_comm_link_i_cast[i].io_clk_tline;
        assign io_valid_tline_li   [i]                       = bsg_comm_link_i_cast[i].io_valid_tline;
        assign io_data_tline_li    [i]                       = bsg_comm_link_i_cast[i].io_data_tline;
        assign bsg_comm_link_o_cast[i].io_token_clk_tline    = io_token_clk_tline_lo[i];
     end

   // out channel
   logic [num_channels_p-1:0]  im_clk_tline_lo;
   logic [num_channels_p-1:0]  im_valid_tline_lo;

   logic [channel_width_p-1:0] im_data_tline_lo [num_channels_p-1:0];
   logic [num_channels_p-1:0]  token_clk_tline_li;

   // output channel conversion
   for (i = 0; i < num_channels_p; i=i+1)
     begin
        assign bsg_comm_link_o_cast[i].im_clk_tline_lo   = im_clk_tline_lo     [i];
        assign bsg_comm_link_o_cast[i].im_valid_tline_lo = im_valid_tline_lo   [i];
        assign bsg_comm_link_o_cast[i].im_data_tline_lo  = im_data_tline_lo    [i];
        assign token_clk_tline_li  [i]                   = bsg_comm_link_i_cast[i].token_clk_tline_li;
     end

   localparam ring_bytes_lp    = 10;
   localparam ring_width_lp = ring_bytes_lp*channel_width_p;

   // **************************************************************
   // *
   // * convert bsg_fsb struct signals to bsg_comm_link format
   // *
   // * fixme: eventually we will push channel grouping down
   // * into bsg_comm_link, but the module is currently in flux
   // *

   `declare_fsb_in_s (ring_width_lp);
   `declare_fsb_out_s(ring_width_lp);

   bsg_fsb_in_s  [nodes_p-1:0] fsb_i_cast;
   bsg_fsb_out_s [nodes_p-1:0] fsb_o_cast;

   assign fsb_i_cast = fsb_i;
   assign fsb_o = fsb_o_cast;

   // into nodes (fsb interface)
   wire [nodes_p-1:0]       core_node_v_A;
   wire [ring_width_lp-1:0] core_node_data_A [nodes_p-1:0];
   wire [nodes_p-1:0]       core_node_ready_A;
    // into nodes (control)
   wire [nodes_p-1:0]      core_node_en_r_lo;
   wire [nodes_p-1:0]      core_node_reset_r_lo;

   // going into nodes (output links of this bsg_comm_link)
   for (i = 0; i < nodes_p; i=i+1)
     begin
        assign fsb_o_cast[i].en_r    = core_node_en_r_lo;
        assign fsb_o_cast[i].reset_r = core_node_reset_r_lo;
        assign fsb_o_cast[i].v       = core_node_v_A   [i];
        assign fsb_o_cast[i].data    = core_node_data_A[i];
        assign core_node_ready_A[i]  = fsb_i_cast[i].ready_rev;
     end

   // out of nodes (input to bsg_comm_link)
   wire [nodes_p-1:0]       core_node_v_B;
   wire [ring_width_lp-1:0] core_node_data_B [nodes_p-1:0];
   wire [nodes_p-1:0]       core_node_yumi_B;

   for (i = 0; i < nodes_p; i=i+1)
     begin
        assign core_node_v_B         [i] = fsb_i_cast[i].v;
        assign core_node_data_B      [i] = fsb_i_cast[i].data;
        assign fsb_o_cast[i].yumi_rev[i] = core_node_ready_B;
     end

   // **************************************************************
   // *
   // * instantiate bsg_comm_link
   // *
   // * fixme: eventually we will push channel grouping down
   // * into bsg_comm_link, but the module is currently in flux
   // *

   // these defaults are appropriate for ASICs, and quick simulation
   // but might be changed for real FPGA or exhaustive simulation

   localparam master_to_slave_speedup_lp = 100;
   localparam snoop_vec_lp               = { nodes_p { 1'b0 } };
   localparam enabled_at_start_vec_lp    = gateway_p;
   localparam master_bypass_test_lp      = 5'b00000;

   bsg_comm_link #(.channel_width_p   (channel_width_p)
                   , .core_channels_p (ring_bytes_lp   )
                   , .link_channels_p (num_channels_p  )
                   , .nodes_p         (nodes_p)
                   , .master_p        (gateway_p)
                   , .master_to_slave_speedup_p(master_to_slave_speedup_lp)
                   , .snoop_vec_p(snoop_vec_lp)
                   , .enabled_at_start_vec_p   (enabled_at_start_vec_lp)
                   , .master_bypass_test_p     (master_bypass_test_lp  )
                   ) comm_link
     (.core_clk_i           (core_clk_i       )
      , .async_reset_i      (async_reset_i    )

      , .io_master_clk_i    (io_master_clk_i  )

      // into nodes (control)
      , .core_node_reset_r_o(core_node_reset_r_lo)
      , .core_node_en_r_o   (core_node_en_r_lo )

      // into nodes (fsb interface)
      , .core_node_v_o      (core_node_v_A    )
      , .core_node_data_o   (core_node_data_A )
      , .core_node_ready_i  (core_node_ready_A)

      // out of nodes (fsb interface)
      , .core_node_v_i   (core_node_v_B   )
      , .core_node_data_i(core_node_data_B)
      , .core_node_yumi_o(core_node_yumi_B)

      // in from i/o
      , .io_valid_tline_i    (io_valid_tline_li    )
      , .io_data_tline_i     (io_data_tline_li     )
      , .io_clk_tline_i      (io_clk_tline_li      )  // clk
      , .io_token_clk_tline_o(io_token_clk_tline_lo)  // clk

      // out to i/o
      , .im_valid_tline_o(im_valid_tline_lo)
      , .im_data_tline_o ( im_data_tline_lo)
      , .im_clk_tline_o  (  im_clk_tline_lo)        // clk

      , .im_slave_reset_tline_r_o (im_slave_reset_tline_r_o)
      , .token_clk_tline_i        (token_clk_tline_li      ) // clk

      ,.core_calib_reset_r_o(core_reset_o)

      // don't use
      , .core_async_reset_danger_o()
      );

endmodule
